// jtag_uart.v

// Generated using ACDS version 13.0sp1 232 at 2025.08.18.22:34:23

`timescale 1 ps / 1 ps
module jtag_uart (
		input  wire        avalon_slave_0_chipselect,  // avalon_slave_0.chipselect
		input  wire        avalon_slave_0_address,     //               .address
		input  wire        avalon_slave_0_read_n,      //               .read_n
		output wire [31:0] avalon_slave_0_readdata,    //               .readdata
		input  wire        avalon_slave_0_write_n,     //               .write_n
		input  wire [31:0] avalon_slave_0_writedata,   //               .writedata
		output wire        avalon_slave_0_waitrequest, //               .waitrequest
		input  wire        clk_in_clk,                 //         clk_in.clk
		input  wire        reset_in_reset              //       reset_in.reset
	);

	jtag_uart_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_in_clk),                 //               clk.clk
		.rst_n          (~reset_in_reset),            //             reset.reset_n
		.av_chipselect  (avalon_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (avalon_slave_0_address),     //                  .address
		.av_read_n      (avalon_slave_0_read_n),      //                  .read_n
		.av_readdata    (avalon_slave_0_readdata),    //                  .readdata
		.av_write_n     (avalon_slave_0_write_n),     //                  .write_n
		.av_writedata   (avalon_slave_0_writedata),   //                  .writedata
		.av_waitrequest (avalon_slave_0_waitrequest), //                  .waitrequest
		.av_irq         ()                            //               irq.irq
	);

endmodule
