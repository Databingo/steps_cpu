// spi.v

// Generated using ACDS version 13.0sp1 232 at 2025.10.10.23:24:13

`timescale 1 ps / 1 ps
module spi (
		input  wire        clk_clk,                           //                    clk.clk
		input  wire        reset_reset_n,                     //                  reset.reset_n
		input  wire        spi_0_reset_reset_n,               //            spi_0_reset.reset_n
		input  wire [15:0] spi_0_spi_control_port_writedata,  // spi_0_spi_control_port.writedata
		output wire [15:0] spi_0_spi_control_port_readdata,   //                       .readdata
		input  wire [2:0]  spi_0_spi_control_port_address,    //                       .address
		input  wire        spi_0_spi_control_port_read_n,     //                       .read_n
		input  wire        spi_0_spi_control_port_chipselect, //                       .chipselect
		input  wire        spi_0_spi_control_port_write_n,    //                       .write_n
		input  wire        spi_0_external_MISO,               //         spi_0_external.MISO
		output wire        spi_0_external_MOSI,               //                       .MOSI
		output wire        spi_0_external_SCLK,               //                       .SCLK
		output wire        spi_0_external_SS_n                //                       .SS_n
	);

	spi_spi_0 spi_0 (
		.clk           (clk_clk),                           //              clk.clk
		.reset_n       (spi_0_reset_reset_n),               //            reset.reset_n
		.data_from_cpu (spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (spi_0_spi_control_port_address),    //                 .address
		.read_n        (spi_0_spi_control_port_read_n),     //                 .read_n
		.spi_select    (spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (spi_0_spi_control_port_write_n),    //                 .write_n
		.irq           (),                                  //              irq.irq
		.MISO          (spi_0_external_MISO),               //         external.export
		.MOSI          (spi_0_external_MOSI),               //                 .export
		.SCLK          (spi_0_external_SCLK),               //                 .export
		.SS_n          (spi_0_external_SS_n)                //                 .export
	);

endmodule
