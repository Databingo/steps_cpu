`define Rom_base  32'h0000_0000
`define Rom_size  32'h0000_0010
`define Ram_base  32'h0000_0010
`define Ram_size  32'h0000_1000
`define Art_base  32'h0000_1010
`define Key_base  32'h0000_1011
