module xhlsTOP
	(
		////////////////////	Clock Input	 	////////////////////	 
		clk27,						//	27 MHz
		RE_N,
		////////////////////	Push Button		////////////////////
		KEY,							//	Pushbutton[5:0]
		////////////////////	DPDT SWitch		////////////////////
		SW,								//	Toggle  SWitch[11:0]
		////////////////////	7-SEG Dispaly	////////////////////
		HEX0,							//	Seven Segment Digit 0
		HEX1,							//	Seven Segment Digit 1
		HEX2,							//	Seven Segment Digit 2
		HEX3,							//	Seven Segment Digit 3
		////////////////////////	LED		////////////////////////
		LEDG,							//	LED Green[7:0]
		LEDR							//	LED Red[11:0]
		////////////////////////	UART	////////////////////////
	);

////////////////////////	Clock Input	 	////////////////////////
input	clk27;				//	27 MHz
input   RE_N;
////////////////////////	Push Button		////////////////////////
input	[5:0]	KEY;					//	Pushbutton[5:0]
////////////////////////	DPDT  SWitch		////////////////////////
input   [11:0]	SW;						//	Toggle  SWitch[11:0]
////////////////////////	7-SEG Dispaly	////////////////////////
output	[6:0]	HEX0;					//	Seven Segment Digit 0
output	[6:0]	HEX1;					//	Seven Segment Digit 1
output	[6:0]	HEX2;					//	Seven Segment Digit 2
output	[6:0]	HEX3;					//	Seven Segment Digit 3
////////////////////////////	LED		////////////////////////////
output	[7:0]	LEDG;					//	LED Green[7:0]
output	[11:0]	LEDR;					//	LED Red[11:0]
///////////////////////////////////////////////////////////////////
wire  [15:0]  mSEG7_DIG;
wire  [15:0]  ouSEG7_DIG;
wire   [7:0]  mtDAA;

wire  [6:0]   mCOUNT;
wire  [7:0]   mDATA;
reg   [23:0]  Cont;

reg       flge;
reg       writ;
reg   [22:0]   Co;
reg   [22:0]   coo;
reg   [22:0]   boo;
reg   [22:0]   goo;
reg   [22:0]   uoo;
reg   [22:0]   doo;
reg   [22:0]   uo;
reg   [22:0]   ddo;
reg   [22:0]   vo;
reg   [22:0]   bo;
reg   [22:0]   eo;
reg   [22:0]   fo;
reg   [22:0]   ffo;
reg   [22:0]   lcdfo;

reg   [22:0]   go;
reg       gkz;
reg       ekz;
reg       fkz;
reg       ffkz;
reg       lcdr;
reg       lcdfkz;

reg       bkz;
reg       kz;     //����ʱ��
reg       vkz;
reg       upkz;
reg       dkz;
reg      bak;
reg      fw;
reg      rest;
reg      clar;
reg      bclar;
reg      lcdclar;

reg      lcdck;

reg      mUP;
reg      mDOWN;
///////////////////////////////////////////////////////////////
assign  LEDR[11]		= SW[0] ? SW[10]  : ouSEG7_DIG[7];
assign  LEDR[10]		= SW[0] ? SW[11]  : ouSEG7_DIG[6];
assign  LEDR[9:4]	   	= SW[0] ? SW[9:4] : ouSEG7_DIG[5:0];
assign  LEDR[3:0]		= SW[3:0];
/*
assign	LEDG[7]	=	~RE_N;
assign	LEDG[6]	=	1'b0;
assign	LEDG[5:0]	=	~KEY[5:0];
//assign	DQ		=	lcdSEG7_DIG;
//assign  gai   = SW[0];*/
assign LEDG[7:0] = mDATA[7:0];

assign	mSEG7_DIG[6]	=  SW[0] ? SW[11]		: ouSEG7_DIG[6];
assign	mSEG7_DIG[7]	=  SW[0] ? SW[10]		: ouSEG7_DIG[7];
assign	mSEG7_DIG[5:0]	=  SW[0] ? SW[9:4]		: ouSEG7_DIG[5:0];
assign	mSEG7_DIG[15]   =  SW[0] ? (SW[1]  ? 1'b0 : mDATA[7]): ouSEG7_DIG[15];
assign	mSEG7_DIG[14:8] =  SW[0] ? ( SW[1] ? mCOUNT[6:0] :	mDATA[6:0])	: ouSEG7_DIG[14:8];


always@(posedge clk18 or negedge RE_N)	
begin
   if (!RE_N)
   begin
     Cont	<=0;
   end
   else
   begin
	  Cont	<=	Cont+1'b1;
      if (mCOUNT!=0)         //����
      begin
	     Cont[23]<=	1'b0;
	     flge <=1'b0;
	  end
      else  flge <=Cont[23];
   end
end

always@(posedge clk18)	
//ȥ����
begin
 
    if (  SW[0]==1 && KEY[2]==0 && kz==0)  //����������
       begin
           Co  <= Co+1'b1;        //���¼�ʱ        
           if (Co==10800 )  writ<=1;
           else  
              begin
                writ <= 0;
                if (Co[22]==1)
                   begin
                    kz<=1;      //ȡֵ��ɱ�־
                    coo<=0;
                   end
              end 
      end 
    else
      begin
         Co<=0;
         writ <= 0;
         coo <= coo+1'b1;
         if (coo[22]==1) kz <= 0;
      end

    if ( SW[0]==1 && KEY[4]==0 && bkz==0)  //�����º���
        begin
           bo<=	bo+1'b1;        //���¼�ʱ        
           if (bo==10800 )   bak<=1;
           else  
              begin
                bak <= 0;
                if ( bo[22]==1'b1 )
                   begin
                    bkz<=1;      //ȡֵ��ɱ�־
                    boo<=0;
                   end
              end 
        end
    else
      begin
         bkz<=1;
         bo<=0;
         bak <= 0;  
         boo <= boo+1'b1;
         if ( boo[22]==1'b1) bkz <= 0;
      end

  if ( SW[0]==1 && KEY[3]==0 && gkz==0)  //������ǰ��
        begin
           go<=	go+1'b1;        //���¼�ʱ        
           if (go==10800)   fw<=1;
           else  
              begin
                fw <= 0;
                if ( go[22]==1'b1 )
                   begin
                    gkz<=1;      //ȡֵ��ɱ�־
                    goo<=0;
                   end
              end 
        end
    else
      begin
         gkz<=1;
         go<=0;
         fw <= 0;  
         goo <= goo+1'b1;
         if ( goo[22]==1'b1) gkz <= 0;
      end
    if ( SW[0]==0  && KEY[4]==0 && upkz==0)  //������ɾ��
        begin
           uo<=	uo+1'b1;        //���¼�ʱ        
           if (uo==10800 )   mUP<=1;
           else  
              begin
                mUP <= 0;
                if ( uo[22]==1'b1 )
                   begin
                    upkz<=1;      //ȡֵ��ɱ�־
                    uoo<=0;
                   end
              end 
        end
    else
      begin
         upkz<=1;
         uo<=0;
         mUP <= 0;  
         uoo <= uoo+1'b1;
         if ( uoo[22]==1'b1) upkz <= 0;
      end

  if ( SW[0]==0  && KEY[3]==0 && dkz==0)  //�����²���
        begin
           ddo<=	ddo+1'b1;        //���¼�ʱ        
           if (ddo==10800 )   mDOWN<=1;
           else  
              begin
                mDOWN <= 0;
                if ( ddo[22]==1'b1 )
                   begin
                    dkz<=1;      //ȡֵ��ɱ�־
                    doo<=0;
                   end
              end 
        end
    else
      begin
         dkz<=1;
         ddo<=0;
         mDOWN <= 0;  
         doo <= doo+1'b1;
         if ( doo[22]==1'b1) dkz <= 0;
      end

    if ( SW[0]==0 && KEY[1]==0)  //������ִ��
        begin
           eo<=	eo+1'b1;        //���¼�ʱ        
           if ((eo==10800 ) && ekz==0) 
              begin
                rest<=1;
                if (eo==10801)
                    ekz<=1; //ȡֵ��־
              end 
              else
                 rest <= 0;
         end
    else
      begin
        ekz<=0;
        eo<=0;
        rest  <= 0;  
      end
    if ( SW[0]==1 && RE_N==0)  //�����¸�λ
        begin
           vo<=	vo+1'b1;        //���¼�ʱ        
           if ((vo==10800  )&& vkz==0) 
              begin
                bclar<=0;
                if (vo==10801)
                vkz<=1; //ȡֵ��־
              end 
              else
                 bclar <= 1;
         end
    else
      begin
        vkz<=0;
        vo<=0;
       bclar  <= 1;  
      end


    if ( SW[0]==0 && RE_N==0)  //�����¸�λ
        begin
           fo<=	fo+1'b1;        //���¼�ʱ        
           if ((fo==10800 )&& fkz==0) 
              begin
                clar<=0;
                if (fo==10801)
                fkz<=1; //ȡֵ��־
              end 
              else
                 clar <= 1;
         end
    else
      begin
        fkz<=0;
        fo<=0;
       clar  <= 1;  
      end

  end 

//����CPU�뻺��������ģ���ʱ�ӣ�
buffcpu  cpu0 (.brak( SW[0]),.clk(clk18),.clr(clar),.wre(writ),
.forw(fw),.back(bak),.data( {SW[10],SW[11],SW[9:4]}),.ol(ouSEG7_DIG[7:0]),
.oh(ouSEG7_DIG[15:8]),.count(mCOUNT),.qb(mDATA));

SEG7_LUT_4 			u0	(	HEX0,HEX1,HEX2,HEX3,mSEG7_DIG,flge);
altpll0 altp0 (.inclk0(clk27),.c0(clk18));


endmodule
