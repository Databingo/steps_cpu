// jtag_uart_system.v

// Generated using ACDS version 13.0sp1 232 at 2025.08.20.23:51:26

`timescale 1 ps / 1 ps
module jtag_uart_system (
		input  wire        clk_clk,                                   //                           clk.clk
		input  wire        reset_reset_n,                             //                         reset.reset_n
		input  wire        jtag_uart_0_avalon_jtag_slave_chipselect,  // jtag_uart_0_avalon_jtag_slave.chipselect
		input  wire        jtag_uart_0_avalon_jtag_slave_address,     //                              .address
		input  wire        jtag_uart_0_avalon_jtag_slave_read_n,      //                              .read_n
		output wire [31:0] jtag_uart_0_avalon_jtag_slave_readdata,    //                              .readdata
		input  wire        jtag_uart_0_avalon_jtag_slave_write_n,     //                              .write_n
		input  wire [31:0] jtag_uart_0_avalon_jtag_slave_writedata,   //                              .writedata
		output wire        jtag_uart_0_avalon_jtag_slave_waitrequest  //                              .waitrequest
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> jtag_uart_0:rst_n

	jtag_uart_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),           //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (jtag_uart_0_avalon_jtag_slave_read_n),      //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (jtag_uart_0_avalon_jtag_slave_write_n),     //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                           //               irq.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
