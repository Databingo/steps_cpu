`define Rom_base  32'h0000_0000
`define Rom_size  32'h0000_0004
`define Ram_base  32'h0000_0004
`define Ram_size  32'h0000_1000
`define Art_base  32'h0000_1004
`define Key_base  32'h0000_1008
