module cpu_on_board (
    (* chip_pin = "PIN_L1" *)  input wire CLOCK_50, // 50 MHz clock
    (* chip_pin = "PIN_R22" *) input wire KEY0,     // Active-low reset button
    (* chip_pin = "PIN_Y21, PIN_Y22, PIN_W21, PIN_W22, PIN_V21, PIN_V22, PIN_U21, PIN_U22" *) output wire [7:0] LEDG, // 8 green LEDs
    (* chip_pin = "R17" *) output reg LEDR9, // 1 red LEDs breath left most 
    (* chip_pin = "U18, Y18, V19, T18, Y19, U19, R19, R20" *) output wire [7:0] LEDR7_0 // 8 red LEDs right
    //(* chip_pin = "R17, R18, U18, Y18, V19, T18, Y19, U19, R19, R20" *) output reg [9:0] LEDR // 10 red LEDs  
);

    (* ram_style = "block" *) reg [31:0] mem [0:2999]; // Unified Memory
    initial $readmemb("mem.mif", mem);

    reg [24:0] counter;
    reg [31:0] addr_pc;
    //
    reg [31:0] ir;
    wire [31:0] ir_bd; assign ir_bd = mem[pc>>2];
    wire [31:0] ir_ld; assign ir_ld = {ir_bd[7:0], ir_bd[15:8], ir_bd[23:16], ir_bd[31:24]};

    reg [31:0] pc;
    reg [63:0] re [0:31]; // General-purpose registers (x0-x31)

    wire clock_1hz;
    clock_slower clock_ins(
	.clk_in(CLOCK_50),
	.clk_out(clock_1hz),
	.reset_n(KEY0)
    );

    // --- Immediate decoders --- 
    wire signed [63:0] w_imm_i = {{52{ir[31]}}, ir[31:20]};   // I-type immediate Lb Lh Lw Lbu Lhu Lwu Ld Jalr Addi Slti Sltiu Xori Ori Andi Addiw
    wire signed [63:0] w_imm_s = {{52{ir[31]}}, ir[31:25], ir[11:7]};  // S-type immediate Sb Sh Sw Sd
    wire signed [63:0] w_imm_b = {{51{ir[31]}}, ir[7],  ir[30:25], ir[11:8], 1'b0}; // SB-type immediate Beq Bne Blt Bge Bltu Bgeu // read immediate & padding last 0, total 12 + 1 = 13 bits
    wire signed [63:0] w_imm_u = {{32{ir[31]}}, ir[31:12], 12'b0}; // U-type immediate Lui Auipc
    wire signed [63:0] w_imm_j = {{43{ir[31]}}, ir[19:12], ir[20], ir[30:21], 1'b0}; // UJ-type immediate Jal  // read immediate & padding last 0, total 20 + 1 = 21 bits
  
    // --- Instruction Decoding ---
    //wire [ 6:0] w_op = ir[6:0];
    wire [ 4:0] w_rd = ir[11:7];
    //wire [ 2:0] w_f3 = ir[14:12]; 
    //wire [ 4:0] w_rs1 = ir[19:15];
    //wire [ 4:0] w_rs2 = ir[24:20];
    //wire [ 6:0] w_f7 = ir[31:25];
    //wire [ 5:0] w_shamt = ir[25:20]; // If 6 bits the highest is always 0??
    //wire [11:0] w_csr = ir[31:20];   // CSR address
    //wire [11:0] w_f12 = ir[31:20];   // ecall 0, ebreak 1
    //wire [ 4:0] w_zimm = ir[19:15];  // CSR zimm

    // IF ir (only fetch)
    always @(posedge clock_1hz or negedge KEY0) begin
        if (!KEY0) begin 
	    LEDR9 <= 1'b0; 
	    ir <= 32'h00000000; 
	end
        else begin
	    LEDR9 <= ~LEDR9; // heartbeat
	    ir <= ir_ld;
        end
    end

    // EXE pc (only one always driver a net)
    always @(posedge clock_1hz or negedge KEY0) begin
        if (!KEY0) begin 
	    pc <=0;
	end
	else begin
	    pc <= pc + 4;
            re[31] <= 1'b0;
    	    casez(ir) 
	    // U-type
            //32'b???????_?????_?????_???_?????_0110111: re[w_rd] <= w_imm_u; // Lui
            //32'b???????_?????_?????_???_?????_0000111: LEDR9 <= 1'b1;
            //32'b???????_?????_?????_???_?????_0110111:  LEDR9 <= 1'b1;
            //32'b???????_?????_?????_???_?????_0110111:  re[0] <= 1'b1;
            //32'b???????_?????_?????_???_?????_0110111:  re[31] <= w_imm_u;
            //32'b???????_?????_?????_???_?????_0110111:  re[31] <= w_rd;
            32'b???????_?????_?????_???_?????_0110111:  re[w_rd] <= w_imm_u;
	    endcase
	end
    end

   assign LEDG = ir[7:0];
   //assign LEDR7_0 = re[31][7:0];
   assign LEDR7_0 = re[31][19:12];



    // Memory controller 
    //always @(posedge clock_1hz or negedge KEY0) begin
    //end

endmodule

<<<<<<< HEAD
=======
// --- TOP ---
module cpu_on_board (
    (* chip_pin = "PIN_L1" *)  input  wire CLOCK_50,
    (* chip_pin = "PIN_R22" *) input  wire KEY0,
    (* chip_pin = "PIN_Y21, PIN_Y22, PIN_W21, PIN_W22, PIN_V21, PIN_V22, PIN_U21, PIN_U22" *)
    output wire [7:0] LEDG,
    (* chip_pin = "R17" *) output wire LEDR9,
    (* chip_pin = "A15" *) output wire TCK,
    (* chip_pin = "B15" *) output wire TMS,
    (* chip_pin = "C15" *) output wire TDI,
    (* chip_pin = "B16" *) output wire TDO
);
    // memory
    (* ram_style = "block" *) reg [31:0] mem [0:2999];
    initial $readmemb("mem.mif", mem);
>>>>>>> 2de6e021648c076659e79e006d9d25c97af50a74



<<<<<<< HEAD

module clock_slower(
    input wire clk_in,
    input wire reset_n,
    output reg clk_out
=======
    // simple “bus”
    reg  [63:0] mem_addr;
    reg  [63:0] mem_data_out;
    reg         mem_we;
    wire [31:0] i_mem_data_in;

    // “UART” write when addr[31]==1
    wire uart_write_en = mem_we && mem_addr[31];

    // NOTE: tck/tms/tdi/tdo are unconnected here; this is a placeholder.
    simple_jtag_uart_tx jtag_uart_inst (
        .tck(TCK), 
	.tms(TMS), 
	.tdi(TDI), 
	.tdo(TDO),   // TODO: replace with a real JTAG/Virtual JTAG
        .clk(CLOCK_50),
        .reset_n(KEY0),
        .write_en(uart_write_en),
        .write_data(mem_data_out[7:0])
>>>>>>> 2de6e021648c076659e79e006d9d25c97af50a74
    );

    reg [24:0] counter; 

    initial begin
	clk_out <= 0;
	counter <=0;
    end

    always @(posedge clk_in or negedge reset_n) begin
	if (!reset_n) begin
	    clk_out <= 0;
	    counter <=0;
	end
	else begin
	    if (counter == 25000000 - 1) begin
		counter <= 0;
		clk_out <= ~clk_out;
	    end
	    else begin
		counter <= counter + 1;
	    end
	end
    end
endmodule



