// =================================================================================
// Original CPU file with minimal changes to force-send 'H' every clock cycle.
// =================================================================================

module cpu_on_board (
    // -- Pin --
    (* chip_pin = "PIN_L1" *)  input wire CLOCK_50, // 50 MHz clock
    (* chip_pin = "PIN_R22" *) input wire KEY0,     // Active-low reset button
    (* chip_pin = "PIN_Y21, PIN_Y22, PIN_W21, PIN_W22, PIN_V21, PIN_V22, PIN_U21, PIN_U22" *) output wire [7:0] LEDG, // 8 green LEDs
    (* chip_pin = "R17" *) output reg LEDR9, // 1 red LEDs breath left most 
    (* chip_pin = "U18, Y18, V19, T18, Y19, U19, R19, R20" *) output wire [7:0] LEDR7_0, // 8 red LEDs right

    (* chip_pin = "H15" *)  input wire PS2_CLK, 
    (* chip_pin = "J14" *)  input wire PS2_DAT 
);

    // -- RAM --
    (* ram_style = "block" *) reg [31:0] mem [0:2999]; // Unified Memory
    initial $readmemb("mem.mif", mem);

    wire [31:0] ir_bd; assign ir_bd = mem[pc>>2];
    wire [31:0] ir_ld; assign ir_ld = {ir_bd[7:0], ir_bd[15:8], ir_bd[23:16], ir_bd[31:24]}; // Endianness swap

riscv64 cpu (
    .clk(clock_1hz), 
    .reset(KEY0),     // Active-low reset button
    .instruction(ir_ld),
    .pc(pc),
    .ir(LEDG),
    //.re(re),
    .heartbeat(LEDR9)
);

   //assign LEDG = ir[7:0];
   //assign LEDR7_0 = re[31][19:12];
   
module riscv64(
    input wire clk, 
    input wire reset,     // Active-low reset button
    input wire [31:0] instruction,
    output reg [31:0] pc,
    output reg [31:0] ir,
    output reg [63:0] re [0:31],
    output wire  heartbeat
);

    
    // --- Immediate decoders (Unchanged) --- 
    wire signed [63:0] w_imm_u = {{32{ir[31]}}, ir[31:12], 12'b0};
    wire [4:0] w_rd  = ir[11:7];

    // IF ir (Unchanged)
    always @(posedge clk or negedge reset) begin
        if (!reset) begin 
            heartbeat <= 1'b0; 
            ir <= 32'h00000000; 
        end else begin
            heartbeat <= ~heartbeat; // heartbeat
            //ir <= ir_ld;
            ir <= instruction;
        end
    end

    // EXE pc (Unchanged, CPU runs normally)
    always @(posedge clk or negedge reset) begin
        if (!reset) begin 
            pc <= 0;
        end else begin
            pc <= pc + 4;
            re[31] <= 1'b0; // This was in your original code
            
	    //data <= 32'h48;
            casez(ir) 
		32'b???????_?????_?????_???_?????_0110111:  re[w_rd] <= w_imm_u; // Lui
		//32'b???????_?????_?????_???_?????_0110111:  begin re[w_rd] <= w_imm_u; data <= 32'h41; end
            endcase
        end
    end

endmodule
   
    // -- Clock --
    wire clock_1hz;
    clock_slower clock_ins(
        .clk_in(CLOCK_50),
        .clk_out(clock_1hz),
        .reset_n(KEY0)
    );

    
   reg [31:0] data;
   wire key_pressed;
   wire key_released;
   reg key_pressed_delay;
   always @(posedge CLOCK_50) begin key_pressed_delay <= key_pressed; end
   ps2_decoder ps2_decoder_inst (
       .clk(CLOCK_50),
       .ps2_clk_async(PS2_CLK),
       .ps2_data_async(PS2_DAT),
       //.scan_code(data[7:0])
       .ascii_code(data[7:0]),
       .key_pressed(key_pressed),
       .key_released(key_released)
   );

    // --- Wires for Avalon-MM Interface (Unchanged from previous JTAG version) ---
    wire [0:0]  avalon_address;
    wire        avalon_write;
    wire [31:0] avalon_writedata;

    // --- Qsys System Instantiation (Unchanged from previous JTAG version) ---
    jtag_uart_system my_jtag_system (
        .clk_clk                             (CLOCK_50),
        .reset_reset_n                       (KEY0),
        .jtag_uart_0_avalon_jtag_slave_address   (avalon_address),
        .jtag_uart_0_avalon_jtag_slave_writedata (avalon_writedata),
        .jtag_uart_0_avalon_jtag_slave_write_n   (~avalon_write),
        .jtag_uart_0_avalon_jtag_slave_chipselect(1'b1),
        .jtag_uart_0_avalon_jtag_slave_read_n    (1'b1)
    );

   wire key_pressed_edge = key_pressed && !key_pressed_delay;
   assign avalon_write     = key_pressed_edge; // Force the write signal high every cycle
   assign avalon_address   = 1'b0;            // Always write to the data register (address 0)
   assign avalon_writedata = {24'b0, data};    

endmodule
