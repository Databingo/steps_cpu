module move_4 (	oSEG0,oSEG1,oSEG2,oSEG3,iDIG,flash,clk );
input	[15:0]	iDIG;		//�����16λ��
input   flash;		//��˸����
input	clk;				//ʱ��
output	[6:0]	oSEG0,oSEG1,oSEG2,oSEG3;	//�����7λ��
reg  [15:0]  dig;
reg  [3:0]  tim;
 
always @(posedge clk)
begin
 dig <= iDIG;
 tim <= tim + 1;
 if (tim[3]) dig <= {dig[11:0],dig[15:12]};
end

SEG7_LUT	u0	(	oSEG0,dig[3:0],flash);		//����һ���������������
SEG7_LUT	u1	(	oSEG1,dig[7:4],flash);
SEG7_LUT	u2	(	oSEG2,dig[11:8],flash);
SEG7_LUT	u3	(	oSEG3,dig[15:12],flash);

endmodule
