module bufuucpu (go,		//�ָ�����
				data,		//��������
				wre,		//дʹ��
				back,		//������
				forw,		//��ǰ���
				clk,		//ʱ��
				clr,		//��λ
				brak,		//�ж�
				oh,			//������ֽ�
				ol,			//������ֽ�
				q,			//�������
				count		//����������
				);
input go,wre,back,forw,clk,clr,brak;
input [7:0] data;
output [7:0] oh,ol,q;
output [6:0] count;
wire w1,w2,w3,w4,w5,irup;		//�м����
wire [7:0] w6;
assign w2=~(brak|irup);  		//�����źŹ�ͬ����

	DFF dff0 (						//����ʱ�괥����
				.d(w1), 			//�������ӣ���֤�ȶ����
				.clk(clk), 
				.clrn(w2), 			//�͵�λ��Ч
				.prn(go), 			//�͵�λ��Ч
				.q(w1)
				);
	//����CPU��			
	jb_cpu cpu0(.clock(clk),.reset_n(clr),.brak(brak),.reset(w1),.read(w3),
		.empty(w4),.orup(irup),.endf(w5),.data(w6),.o({oh,ol}));
//���û�������
	buffin buff0(.data(data),.wre(wre),.back(back),.clk(clk),.clr(clr),
		.read(w3),.forw(forw),.empt(w4),.endf(w5),.q(q),.count(count),
		.out(w6));
endmodule 
