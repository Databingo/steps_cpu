`define Rom_base  32'h0000_0000
`define Rom_size  32'h0000_1000; // 4KB ROM
`define Ram_base  32'h0000_1000
`define Ram_size  32'h0000_2000; // 4KB RAM
`define Art_base  32'h0000_ffff; 
`define Key_base  32'h0000_fffe; 
