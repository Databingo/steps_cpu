// sd.v

// Generated using ACDS version 13.0sp1 232 at 2025.10.15.01:54:39

`timescale 1 ps / 1 ps
module sd (
		input  wire        clk_clk,                                                              //                                                      clk.clk
		input  wire        reset_reset_n,                                                        //                                                    reset.reset_n
		inout  wire        altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_cmd,            //         altera_up_sd_card_avalon_interface_0_conduit_end.b_SD_cmd
		inout  wire        altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat,            //                                                         .b_SD_dat
		inout  wire        altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat3,           //                                                         .b_SD_dat3
		output wire        altera_up_sd_card_avalon_interface_0_conduit_end_o_SD_clock,          //                                                         .o_SD_clock
		input  wire        altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,  // altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave.chipselect
		input  wire [7:0]  altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,     //                                                         .address
		input  wire        altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,        //                                                         .read
		input  wire        altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,       //                                                         .write
		input  wire [3:0]  altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,  //                                                         .byteenable
		input  wire [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,   //                                                         .writedata
		output wire [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,    //                                                         .readdata
		output wire        altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest  //                                                         .waitrequest
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (clk_clk),                                                              //          clock_sink.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                                      //    clock_sink_reset.reset_n
		.b_SD_cmd             (altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_cmd),            //         conduit_end.export
		.b_SD_dat             (altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat),            //                    .export
		.b_SD_dat3            (altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat3),           //                    .export
		.o_SD_clock           (altera_up_sd_card_avalon_interface_0_conduit_end_o_SD_clock)           //                    .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
